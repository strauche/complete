dut.v