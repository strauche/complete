package tests_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import env_pkg::*;
  import my_pkg::*;

  `include "my_test.sv"
  `include "test1.sv"
  `include "test2.sv"
  `include "test3.sv"

endpackage: tests_pkg
